* C:\Users\kumar\eSim-Workspace\double_tail_comp\double_tail_comp.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/09/22 16:01:43

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  outp Net-_M1-Pad2_ GND GND mosfet_n		
M5  outp outn GND GND mosfet_n		
M8  outn outp GND GND mosfet_n		
M12  outn Net-_M10-Pad1_ GND GND mosfet_n		
M3  outp outn Net-_M11-Pad3_ Net-_M11-Pad3_ mosfet_p		
M11  outn outp Net-_M11-Pad3_ Net-_M11-Pad3_ mosfet_p		
M7  Net-_M11-Pad3_ Net-_M7-Pad2_ vdd vdd mosfet_p		
M2  Net-_M1-Pad2_ clk vdd vdd mosfet_p		
M10  Net-_M10-Pad1_ clk vdd vdd mosfet_p		
M4  Net-_M1-Pad2_ in1 Net-_M4-Pad3_ GND mosfet_n		
M9  Net-_M10-Pad1_ in2 Net-_M4-Pad3_ GND mosfet_n		
M6  Net-_M4-Pad3_ clk GND GND mosfet_n		
v1  clk GND pulse		
v2  vdd GND 5		
v4  in1 GND sine		
X1  clk Net-_M7-Pad2_ INVCMOS		
v3  in2 GND 1		

.end
