* C:\Users\kumar\eSim-Workspace\dtc__new\dtc__new.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/10/22 21:38:23

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  vref vr1 10k		
R2  vr1 vr2 10k		
R3  vr2 vr3 10k		
R4  vr3 vr4 10k		
R5  vr4 vr5 10k		
R6  vr5 vr6 10k		
R7  vr6 vr7 10k		
R8  vr7 GND 10k		
v2  vdd GND 14		
v3  vref GND 1		
v1  vin GND sine		
X5  ? vr1 vin vss ? o1 vdd ? lm_741		
X6  ? vr2 vin vss ? o2 vdd ? lm_741		
X2  ? vr3 vin vss ? o3 vdd ? lm_741		
X3  ? vr4 vin vss ? o4 vdd ? lm_741		
X4  ? vr5 vin vss ? o5 vdd ? lm_741		
X1  ? vr7 vin vss ? o7 vdd ? lm_741		
v4  GND vss 14		
X7  ? vr6 vin vss ? o6 vdd ? lm_741		
U5  out1 plot_v1		
U6  out2 plot_v1		
U7  out3 plot_v1		
U2  Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ out1 out2 out3 dac_bridge_3		
U3  o1 o2 o3 o4 o5 o6 o7 GND Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ adc_bridge_8		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ charaan_pe		

.end
